`timescale 1ns / 1ps

module convolverlayer2(clk,ce,weight1,global_rst,activation1,bias,end_activate,data_out,valid_conv,outcount1,maxout);
//parameter n = 32'd512;     // activation map size->input size
parameter k = 9'd3;     // kernel size 
parameter step1 =4'd2;
parameter outlenper=13'd30;
parameter outlenall=13'd1260;
//parameter batch=6'd42;

input wire clk,ce,global_rst;
input wire  [16:0] activation1;
input wire signed   [7:0] bias ;
input wire   [8*k-1:0]weight1;
//output wire [8*outlen-1:0] data_out1;
output wire end_activate;
output wire [31:0] data_out;
output wire valid_conv;
output wire [10:0] outcount1;
output wire [31:0] maxout;
//output wire dataout_begin;
//test pin
//output wire [15:0] conv_op;
//wire clk8;
///////////////////////////////////////////�޸�
//reg [7:0] data_out[0:outlen-1];
reg signed [31:0]  data_outreg;
//test
reg  signed [31:0]  maxoutreg;
wire signed [31:0] tmp [0:k];

//reg dataout_beginreg;

wire signed [31:0] conv_op;
//wire [23:0] relu_op;
reg end_activatetem;
assign tmp[0]=0;




assign data_out=data_outreg;
assign maxout=maxoutreg;



generate
genvar i;
for(i = 0;i<k;i=i+1)
begin: MAC
//(* use_dsp = "yes" *)               //this line is optional depending on tool behaviour
MAClayer2 mac2(                     //implements a*b+c
  .clk(clk), // input clk
  .ce(ce), // input ce
  .sclr(global_rst), // input sclr
  .a(activation1), // activation input [15 : 0] a
  .b(weight1[8*i +: 8]), // weight input [15 : 0] b
  .c(tmp[i]), // previous mac sum input [31 : 0] c
  .p(tmp[i+1]) // output [31 : 0] p
  );
end 
//end 
endgenerate

reg [31:0] countclk;
reg [10:0] outcount;
reg [11:0] countper;
//reg [5:0]  outcountbatch;
reg en2,en3;
reg [5:0] step;

assign outcount1=outcount;

integer d;
always@(posedge clk ) begin
if(global_rst)
begin
countclk<=32'b0;     
//countstep<=32'b0;
outcount<=11'b0;
countper<=0;
step<=step1;
//dataout_beginreg<=0;
en2<=1'b0;
en3<=1'b0;
//for(d=0;d<outlen;d=d+1) begin
data_outreg<=0;//end
end_activatetem<=0;
maxoutreg<=0;
end

else if(ce)
    if((countclk>=k-1)) 
//����ʱ�����⣬��һ�������ڵ�K+1�����ڳ��������Ǽ�������һ�����ڣ���Ҫ��ǰһ������Ԥ��en2��poseclkһ��������en3ʧЧ
        begin
            en2 <= 1'b1;
            countclk<= countclk+1'b1;
        end
    else
        begin 
        en2<= 1'b0;
        countclk<= countclk+1'b1;
        end
end

always @(posedge clk)begin
if(global_rst)
outcount<=0;

else begin

if((en2==1))  begin
    if (countclk==k+countper*(k-step)+outcount*step)
        begin
            en3 <= 1'b1;
            if(outcount==outlenall)
           outcount<=outcount;
            else 
            outcount<=outcount+1;
        end
                
/////////////////////////////////////////////////////////////16:46mod
//else if (countclk!=k+1+outcount*step)
    else
           en3<=1'b0;
                    end
 else begin
         outcount<=0;
        en3<=0; 
        end
        end
end
//end
///////////////////////////////


assign valid_conv = (en2&&en3);
assign conv_op=valid_conv?(tmp[k]+bias):0;
//assign end_conv = (count>= n+k)?1'b1:1'b0;

// relu act(valid_conv,conv_op,relu_op);


always@(negedge clk) begin//��Ϊ�½���
  if(valid_conv) 
  begin
//data_out[outcount-1]<={relu_op[15:8]};//����ʱ�������ڵ�120��outcount�Ѿ���1
data_outreg<=conv_op;

////////////test
if(maxoutreg<data_outreg)
maxoutreg<=data_outreg;
 

    if(outcount==outlenper*(countper+1))begin
  //step<=k;
  countper<=countper+1;
  //end_activatetem<=1'b1;
  end
   if(outcount==outlenall)begin
   end_activatetem<=1'b1;end
  
  
  end
end
assign end_activate=end_activatetem;

endmodule
